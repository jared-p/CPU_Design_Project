library verilog;
use verilog.vl_types.all;
entity test_memory_read is
end test_memory_read;
