library verilog;
use verilog.vl_types.all;
entity Test_Registry_Bank is
end Test_Registry_Bank;
