library verilog;
use verilog.vl_types.all;
entity memory_control_with_RAM_testbench is
end memory_control_with_RAM_testbench;
