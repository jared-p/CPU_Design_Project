library verilog;
use verilog.vl_types.all;
entity final_design_test is
end final_design_test;
