library verilog;
use verilog.vl_types.all;
entity Test_ALU is
end Test_ALU;
